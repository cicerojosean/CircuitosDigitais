library verilog;
use verilog.vl_types.all;
entity cronometro_vlg_vec_tst is
end cronometro_vlg_vec_tst;
