library verilog;
use verilog.vl_types.all;
entity horario_vlg_vec_tst is
end horario_vlg_vec_tst;
